module test();



endmodule