module sevenseg (x,s);
	
	input [3:0]x;
	output [6:0]s;	

	assign s[0] = (~x[3] & ~x[2] & ~x[1] & x[0])|(~x[3] & x[2] & ~x[1] & ~x[0])|(x[3] & ~x[2] & x[1] & x[0])|(x[3] & x[2] & ~x[1] & x[0]);
	assign s[1] = (~x[3] & x[2] & ~x[1] & x[0])|(~x[3] & x[2] & x[1] & ~x[0])|(x[3] & ~x[2] & x[1] & x[0])|(x[3] & x[2] & ~x[1] & ~x[0])|(x[3] & x[2] & x[1] & ~x[0])|(x[3] & x[2] & x[1] & x[0]);
	assign s[2] = (~x[3] & ~x[2] & x[1] & ~x[0])|(x[3] & x[2] & ~x[1] & ~x[0])|(x[3] & x[2] & x[1] & ~x[0])|(x[3] & x[2] & x[1] & x[0]);
	assign s[3] = (~x[3] & ~x[2] & ~x[1] & x[0])|(~x[3] & x[2] & ~x[1] & ~x[0])|(~x[3] & x[2] & x[1] & x[0])|(x[3] & ~x[2] & x[1] & ~x[0])|(x[3] & x[2] & x[1] & x[0]);
	assign s[4] = (~x[3] & ~x[2] & ~x[1] & x[0])|(~x[3] & ~x[2] & x[1] & x[0])|(~x[3] & x[2] & ~x[1] & ~x[0])|(~x[3] & x[2] & ~x[1] & x[0])|(~x[3] & x[2] & x[1] & x[0])|(x[3] & ~x[2] & ~x[1] & x[0]);
	assign s[5] = (~x[3] & ~x[2] & ~x[1] & x[0])|(~x[3] & ~x[2] & x[1] & ~x[0])|(~x[3] & ~x[2] & x[1] & x[0])|(~x[3] & x[2] & x[1] & x[0])|(x[3] & x[2] & ~x[1] & x[0]);
	assign s[6] = (~x[3] & ~x[2] & ~x[1])|(~x[3] & ~x[2] & ~x[1])|(~x[3] & x[2] & x[1] & x[0])|(x[3] & x[2] & ~x[1] & ~x[0]);

endmodule