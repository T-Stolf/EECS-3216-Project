module displayLines();// input clock 25MHz horizontal space: 640px (144-783) vertical space: 480px (35-514)

endmodule